`include "mux2to1.v"

module Lshift16(A, shl, OUT);

	input [15:0] A;
	input [3:0] shl;

	output [15:0] OUT;

	wire [15:0] m0, m1, m2, m3;

	reg z = 1'b0;

	mux2to1 M00(z, A[0], ~shl[0], m0[0]), M01(A[0], A[1], ~shl[0], m0[1]), M02(A[1], A[2], ~shl[0], m0[2]), M03(A[2], A[3], ~shl[0], m0[3]), M04(A[3], A[4], ~shl[0], m0[4]), M05(A[4], A[5], ~shl[0], m0[5]), M06(A[5], A[6], ~shl[0], m0[6]), M07(A[6], A[7], ~shl[0], m0[7]), M08(A[7], A[8], ~shl[0], m0[8]), M09(A[8], A[9], ~shl[0], m0[9]), M010(A[9], A[10], ~shl[0], m0[10]), M011(A[10], A[11], ~shl[0], m0[11]), M012(A[11], A[12], ~shl[0], m0[12]), M013(A[12], A[13], ~shl[0], m0[13]), M014(A[13], A[14], ~shl[0], m0[14]), M015(A[14], A[15], ~shl[0], m0[15]);

	mux2to1 M10(z, m0[0], ~shl[1], m1[0]), M11(z, m0[1], ~shl[1], m1[1]), M12(m0[0], m0[2], ~shl[1], m1[2]), M13(m0[1], m0[3], ~shl[1], m1[3]), M14(m0[2], m0[4], ~shl[1], m1[4]), M15(m0[3], m0[5], ~shl[1], m1[5]), M16(m0[4], m0[6], ~shl[1], m1[6]), M17(m0[5], m0[7], ~shl[1], m1[7]), M18(m0[6], m0[8], ~shl[1], m1[8]), M19(m0[7], m0[9], ~shl[1], m1[9]), M110(m0[8], m0[10], ~shl[1], m1[10]), M111(m0[9], m0[11], ~shl[1], m1[11]), M112(m0[10], m0[12], ~shl[1], m1[12]), M113(m0[11], m0[13], ~shl[1], m1[13]), M114(m0[12], m0[14], ~shl[1], m1[14]), M115(m0[13], m0[15], ~shl[1], m1[15]);

	mux2to1 M20(z, m1[0], ~shl[2], m2[0]), M21(z, m1[1], ~shl[2], m2[1]), M22(z, m1[2], ~shl[2], m2[2]), M23(z, m1[3], ~shl[2], m2[3]), M24(m1[0], m1[4], ~shl[2], m2[4]), M25(m1[1], m1[5], ~shl[2], m2[5]), M26(m1[2], m1[6], ~shl[2], m2[6]), M27(m1[3], m1[7], ~shl[2], m2[7]), M28(m1[4], m1[8], ~shl[2], m2[8]), M29(m1[5], m1[9], ~shl[2], m2[9]), M210(m1[6], m1[10], ~shl[2], m2[10]), M211(m1[7], m1[11], ~shl[2], m2[11]), M212(m1[8], m1[12], ~shl[2], m2[12]), M213(m1[9], m1[13], ~shl[2], m2[13]), M214(m1[10], m1[14], ~shl[2], m2[14]), M215(m1[11], m1[15], ~shl[2], m2[15]);

	mux2to1 M30(z, m2[0], ~shl[3], m3[0]), M31(z, m2[1], ~shl[3], m3[1]), M32(z, m2[2], ~shl[3], m3[2]), M33(z, m2[3], ~shl[3], m3[3]), M34(z, m2[4], ~shl[3], m3[4]), M35(z, m2[5], ~shl[3], m3[5]), M36(z, m2[6], ~shl[3], m3[6]), M37(z, m2[7], ~shl[3], m3[7]), M38(m2[0], m2[8], ~shl[3], m3[8]), M39(m2[1], m2[9], ~shl[3], m3[9]), M310(m2[2], m2[10], ~shl[3], m3[10]), M311(m2[3], m2[11], ~shl[3], m3[11]), M312(m2[4], m2[12], ~shl[3], m3[12]), M313(m2[5], m2[13], ~shl[3], m3[13]), M314(m2[6], m2[14], ~shl[3], m3[14]), M315(m2[7], m2[15], ~shl[3], m3[15]);

	assign OUT = m3;

endmodule
