`include "Prefix_Add16.v"

module mult16(x, y, P);

	input [15:0] x, y;

	output [31:0] P;

	reg zero = 1'b0;

	wire [15:0] p0;
	wire [16:1] p1;
	wire [17:2] p2;
	wire [18:3] p3;
	wire [19:4] p4;
	wire [20:5] p5;
	wire [21:6] p6;
	wire [22:7] p7;
	wire [23:8] p8;
	wire [24:9] p9;
	wire [25:10] p10;
	wire [26:11] p11;
	wire [27:12] p12;
	wire [28:13] p13;
	wire [29:14] p14;
	wire [30:15] p15;

	wire [16:0] s0;
	wire [17:1] s1;
	wire [18:2] s2;
	wire [19:3] s3;
	wire [20:4] s4;
	wire [21:5] s5;
	wire [22:6] s6;
	wire [23:7] s7;
	wire [24:8] s8;
	wire [25:9] s9;
	wire [26:10] s10;
	wire [27:11] s11;
	wire [28:12] s12;
	wire [29:13] s13;
	wire [30:14] s14;
	wire [31:15] s15;

	assign s0[16] = zero;

	assign p0[15] = y[0]&x[15], p0[14] = y[0]&x[14], p0[13] = y[0]&x[13], p0[12] = y[0]&x[12], p0[11] = y[0]&x[11], p0[10] = y[0]&x[10], p0[9] = y[0]&x[9], p0[8] = y[0]&x[8], p0[7] = y[0]&x[7], p0[6] = y[0]&x[6], p0[5] = y[0]&x[5], p0[4] = y[0]&x[4], p0[3] = y[0]&x[3], p0[2] = y[0]&x[2], p0[1] = y[0]&x[1], p0[0] = y[0]&x[0];
	assign p1[16] = y[1]&x[15], p1[15] = y[1]&x[14], p1[14] = y[1]&x[13], p1[13] = y[1]&x[12], p1[12] = y[1]&x[11], p1[11] = y[1]&x[10], p1[10] = y[1]&x[9], p1[9] = y[1]&x[8], p1[8] = y[1]&x[7], p1[7] = y[1]&x[6], p1[6] = y[1]&x[5], p1[5] = y[1]&x[4], p1[4] = y[1]&x[3], p1[3] = y[1]&x[2], p1[2] = y[1]&x[1], p1[1] = y[1]&x[0];
	assign p2[17] = y[2]&x[15], p2[16] = y[2]&x[14], p2[15] = y[2]&x[13], p2[14] = y[2]&x[12], p2[13] = y[2]&x[11], p2[12] = y[2]&x[10], p2[11] = y[2]&x[9], p2[10] = y[2]&x[8], p2[9] = y[2]&x[7], p2[8] = y[2]&x[6], p2[7] = y[2]&x[5], p2[6] = y[2]&x[4], p2[5] = y[2]&x[3], p2[4] = y[2]&x[2], p2[3] = y[2]&x[1], p2[2] = y[2]&x[0];
	assign p3[18] = y[3]&x[15], p3[17] = y[3]&x[14], p3[16] = y[3]&x[13], p3[15] = y[3]&x[12], p3[14] = y[3]&x[11], p3[13] = y[3]&x[10], p3[12] = y[3]&x[9], p3[11] = y[3]&x[8], p3[10] = y[3]&x[7], p3[9] = y[3]&x[6], p3[8] = y[3]&x[5], p3[7] = y[3]&x[4], p3[6] = y[3]&x[3], p3[5] = y[3]&x[2], p3[4] = y[3]&x[1], p3[3] = y[3]&x[0];
	assign p4[19] = y[4]&x[15], p4[18] = y[4]&x[14], p4[17] = y[4]&x[13], p4[16] = y[4]&x[12], p4[15] = y[4]&x[11], p4[14] = y[4]&x[10], p4[13] = y[4]&x[9], p4[12] = y[4]&x[8], p4[11] = y[4]&x[7], p4[10] = y[4]&x[6], p4[9] = y[4]&x[5], p4[8] = y[4]&x[4], p4[7] = y[4]&x[3], p4[6] = y[4]&x[2], p4[5] = y[4]&x[1], p4[4] = y[4]&x[0];
	assign p5[20] = y[5]&x[15], p5[19] = y[5]&x[14], p5[18] = y[5]&x[13], p5[17] = y[5]&x[12], p5[16] = y[5]&x[11], p5[15] = y[5]&x[10], p5[14] = y[5]&x[9], p5[13] = y[5]&x[8], p5[12] = y[5]&x[7], p5[11] = y[5]&x[6], p5[10] = y[5]&x[5], p5[9] = y[5]&x[4], p5[8] = y[5]&x[3], p5[7] = y[5]&x[2], p5[6] = y[5]&x[1], p5[5] = y[5]&x[0];
	assign p6[21] = y[6]&x[15], p6[20] = y[6]&x[14], p6[19] = y[6]&x[13], p6[18] = y[6]&x[12], p6[17] = y[6]&x[11], p6[16] = y[6]&x[10], p6[15] = y[6]&x[9], p6[14] = y[6]&x[8], p6[13] = y[6]&x[7], p6[12] = y[6]&x[6], p6[11] = y[6]&x[5], p6[10] = y[6]&x[4], p6[9] = y[6]&x[3], p6[8] = y[6]&x[2], p6[7] = y[6]&x[1], p6[6] = y[6]&x[0];
	assign p7[22] = y[7]&x[15], p7[21] = y[7]&x[14], p7[20] = y[7]&x[13], p7[19] = y[7]&x[12], p7[18] = y[7]&x[11], p7[17] = y[7]&x[10], p7[16] = y[7]&x[9], p7[15] = y[7]&x[8], p7[14] = y[7]&x[7], p7[13] = y[7]&x[6], p7[12] = y[7]&x[5], p7[11] = y[7]&x[4], p7[10] = y[7]&x[3], p7[9] = y[7]&x[2], p7[8] = y[7]&x[1], p7[7] = y[7]&x[0];
	assign p8[23] = y[8]&x[15], p8[22] = y[8]&x[14], p8[21] = y[8]&x[13], p8[20] = y[8]&x[12], p8[19] = y[8]&x[11], p8[18] = y[8]&x[10], p8[17] = y[8]&x[9], p8[16] = y[8]&x[8], p8[15] = y[8]&x[7], p8[14] = y[8]&x[6], p8[13] = y[8]&x[5], p8[12] = y[8]&x[4], p8[11] = y[8]&x[3], p8[10] = y[8]&x[2], p8[9] = y[8]&x[1], p8[8] = y[8]&x[0];
	assign p9[24] = y[9]&x[15], p9[23] = y[9]&x[14], p9[22] = y[9]&x[13], p9[21] = y[9]&x[12], p9[20] = y[9]&x[11], p9[19] = y[9]&x[10], p9[18] = y[9]&x[9], p9[17] = y[9]&x[8], p9[16] = y[9]&x[7], p9[15] = y[9]&x[6], p9[14] = y[9]&x[5], p9[13] = y[9]&x[4], p9[12] = y[9]&x[3], p9[11] = y[9]&x[2], p9[10] = y[9]&x[1], p9[9] = y[9]&x[0];
	assign p10[25] = y[10]&x[15], p10[24] = y[10]&x[14], p10[23] = y[10]&x[13], p10[22] = y[10]&x[12], p10[21] = y[10]&x[11], p10[20] = y[10]&x[10], p10[19] = y[10]&x[9], p10[18] = y[10]&x[8], p10[17] = y[10]&x[7], p10[16] = y[10]&x[6], p10[15] = y[10]&x[5], p10[14] = y[10]&x[4], p10[13] = y[10]&x[3], p10[12] = y[10]&x[2], p10[11] = y[10]&x[1], p10[10] = y[10]&x[0];
	assign p11[26] = y[11]&x[15], p11[25] = y[11]&x[14], p11[24] = y[11]&x[13], p11[23] = y[11]&x[12], p11[22] = y[11]&x[11], p11[21] = y[11]&x[10], p11[20] = y[11]&x[9], p11[19] = y[11]&x[8], p11[18] = y[11]&x[7], p11[17] = y[11]&x[6], p11[16] = y[11]&x[5], p11[15] = y[11]&x[4], p11[14] = y[11]&x[3], p11[13] = y[11]&x[2], p11[12] = y[11]&x[1], p11[11] = y[11]&x[0];
	assign p12[27] = y[12]&x[15], p12[26] = y[12]&x[14], p12[25] = y[12]&x[13], p12[24] = y[12]&x[12], p12[23] = y[12]&x[11], p12[22] = y[12]&x[10], p12[21] = y[12]&x[9], p12[20] = y[12]&x[8], p12[19] = y[12]&x[7], p12[18] = y[12]&x[6], p12[17] = y[12]&x[5], p12[16] = y[12]&x[4], p12[15] = y[12]&x[3], p12[14] = y[12]&x[2], p12[13] = y[12]&x[1], p12[12] = y[12]&x[0];
	assign p13[28] = y[13]&x[15], p13[27] = y[13]&x[14], p13[26] = y[13]&x[13], p13[25] = y[13]&x[12], p13[24] = y[13]&x[11], p13[23] = y[13]&x[10], p13[22] = y[13]&x[9], p13[21] = y[13]&x[8], p13[20] = y[13]&x[7], p13[19] = y[13]&x[6], p13[18] = y[13]&x[5], p13[17] = y[13]&x[4], p13[16] = y[13]&x[3], p13[15] = y[13]&x[2], p13[14] = y[13]&x[1], p13[13] = y[13]&x[0];
	assign p14[29] = y[14]&x[15], p14[28] = y[14]&x[14], p14[27] = y[14]&x[13], p14[26] = y[14]&x[12], p14[25] = y[14]&x[11], p14[24] = y[14]&x[10], p14[23] = y[14]&x[9], p14[22] = y[14]&x[8], p14[21] = y[14]&x[7], p14[20] = y[14]&x[6], p14[19] = y[14]&x[5], p14[18] = y[14]&x[4], p14[17] = y[14]&x[3], p14[16] = y[14]&x[2], p14[15] = y[14]&x[1], p14[14] = y[14]&x[0];
	assign p15[30] = y[15]&x[15], p15[29] = y[15]&x[14], p15[28] = y[15]&x[13], p15[27] = y[15]&x[12], p15[26] = y[15]&x[11], p15[25] = y[15]&x[10], p15[24] = y[15]&x[9], p15[23] = y[15]&x[8], p15[22] = y[15]&x[7], p15[21] = y[15]&x[6], p15[20] = y[15]&x[5], p15[19] = y[15]&x[4], p15[18] = y[15]&x[3], p15[17] = y[15]&x[2], p15[16] = y[15]&x[1], p15[15] = y[15]&x[0];


	assign s0[15:0] = p0;

	Prefix_Add16 f1(s0[16:1], p1[16:1], zero, s1[16:1], s1[17]);
	Prefix_Add16 f2(s1[17:2], p2[17:2], zero, s2[17:2], s2[18]);
	Prefix_Add16 f3(s2[18:3], p3[18:3], zero, s3[18:3], s3[19]);
	Prefix_Add16 f4(s3[19:4], p4[19:4], zero, s4[19:4], s4[20]);
	Prefix_Add16 f5(s4[20:5], p5[20:5], zero, s5[20:5], s5[21]);
	Prefix_Add16 f6(s5[21:6], p6[21:6], zero, s6[21:6], s6[22]);
	Prefix_Add16 f7(s6[22:7], p7[22:7], zero, s7[22:7], s7[23]);
	Prefix_Add16 f8(s7[23:8], p8[23:8], zero, s8[23:8], s8[24]);
	Prefix_Add16 f9(s8[24:9], p9[24:9], zero, s9[24:9], s9[25]);
	Prefix_Add16 f10(s9[25:10], p10[25:10], zero, s10[25:10], s10[26]);
	Prefix_Add16 f11(s10[26:11], p11[26:11], zero, s11[26:11], s11[27]);
	Prefix_Add16 f12(s11[27:12], p12[27:12], zero, s12[27:12], s12[28]);
	Prefix_Add16 f13(s12[28:13], p13[28:13], zero, s13[28:13], s13[29]);
	Prefix_Add16 f14(s13[29:14], p14[29:14], zero, s14[29:14], s14[30]);
	Prefix_Add16 f15(s14[30:15], p15[30:15], zero, s15[30:15], s15[31]);


	assign P[0] = s0[0];
	assign P[1] = s1[1];
	assign P[2] = s2[2];
	assign P[3] = s3[3];
	assign P[4] = s4[4];
	assign P[5] = s5[5];
	assign P[6] = s6[6];
	assign P[7] = s7[7];
	assign P[8] = s8[8];
	assign P[9] = s9[9];
	assign P[10] = s10[10];
	assign P[11] = s11[11];
	assign P[12] = s12[12];
	assign P[13] = s13[13];
	assign P[14] = s14[14];

	assign P[31:15] = s15[31:15];


endmodule
