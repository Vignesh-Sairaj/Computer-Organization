module PC(inout addr);

    
endmodule
