module Prefix_Add8(x, y, cIn, s, cOut);

	input [7:0] x, y;
	input cIn;

	output [7:0] s;
	output cOut;

	wire [7:0] g0, p0, g1, p1, g2, p2, g3, p3;
	wire [8:0] c;

	assign g0[7:1] = x[7:1]&y[7:1];
	assign p0[7:0] = x^y;
	assign c[0] = cIn;
	assign g0[0] = x[0]&y[0] | c[0]&(x[0] | y[0]);



	assign g1[7] = g0[7] | p0[7]&g0[6], g1[6] = g0[6] | p0[6]&g0[5], g1[5] = g0[5] | p0[5]&g0[4], g1[4] = g0[4] | p0[4]&g0[3], g1[3] = g0[3] | p0[3]&g0[2], g1[2] = g0[2] | p0[2]&g0[1], g1[1] = g0[1] | p0[1]&g0[0], g1[0] = g0[0];
	assign p1[7] = p0[7]&p0[6], p1[6] = p0[6]&p0[5], p1[5] = p0[5]&p0[4], p1[4] = p0[4]&p0[3], p1[3] = p0[3]&p0[2], p1[2] = p0[2]&p0[1], p1[1] = p0[1]&p0[0], p1[0] = p0[0];

	assign g2[7] = g1[7] | p1[7]&g1[5], g2[6] = g1[6] | p1[6]&g1[4], g2[5] = g1[5] | p1[5]&g1[3], g2[4] = g1[4] | p1[4]&g1[2], g2[3] = g1[3] | p1[3]&g1[1], g2[2] = g1[2] | p1[2]&g1[0], g2[1] = g1[1], g2[0] = g1[0];
	assign p2[7] = p1[7]&p1[5], p2[6] = p1[6]&p1[4], p2[5] = p1[5]&p1[3], p2[4] = p1[4]&p1[2], p2[3] = p1[3]&p1[1], p2[2] = p1[2]&p1[0], p2[1] = p1[1], p2[0] = p1[0];

	assign g3[7] = g2[7] | p2[7]&g2[3], g3[6] = g2[6] | p2[6]&g2[2], g3[5] = g2[5] | p2[5]&g2[1], g3[4] = g2[4] | p2[4]&g2[0], g3[3] = g2[3], g3[2] = g2[2], g3[1] = g2[1], g3[0] = g2[0];
	assign p3[7] = p2[7]&p2[3], p3[6] = p2[6]&p2[2], p3[5] = p2[5]&p2[1], p3[4] = p2[4]&p2[0], p3[3] = p2[3], p3[2] = p2[2], p3[1] = p2[1], p3[0] = p2[0];



	assign c[8:1] = g3[7:0];
	assign s = p0^c[7:0];
	assign cOut = c[8];

endmodule
