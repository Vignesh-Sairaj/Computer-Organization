`include "Prefix_Add32.v"

module Array_Mult32_gen(x, y, P);

	input [31:0] x, y;

	output [63:0] P;

	reg zero = 1'b0;

	wire [31:0] p0;
	wire [32:1] p1;
	wire [33:2] p2;
	wire [34:3] p3;
	wire [35:4] p4;
	wire [36:5] p5;
	wire [37:6] p6;
	wire [38:7] p7;
	wire [39:8] p8;
	wire [40:9] p9;
	wire [41:10] p10;
	wire [42:11] p11;
	wire [43:12] p12;
	wire [44:13] p13;
	wire [45:14] p14;
	wire [46:15] p15;
	wire [47:16] p16;
	wire [48:17] p17;
	wire [49:18] p18;
	wire [50:19] p19;
	wire [51:20] p20;
	wire [52:21] p21;
	wire [53:22] p22;
	wire [54:23] p23;
	wire [55:24] p24;
	wire [56:25] p25;
	wire [57:26] p26;
	wire [58:27] p27;
	wire [59:28] p28;
	wire [60:29] p29;
	wire [61:30] p30;
	wire [62:31] p31;

	wire [32:0] s0;
	wire [33:1] s1;
	wire [34:2] s2;
	wire [35:3] s3;
	wire [36:4] s4;
	wire [37:5] s5;
	wire [38:6] s6;
	wire [39:7] s7;
	wire [40:8] s8;
	wire [41:9] s9;
	wire [42:10] s10;
	wire [43:11] s11;
	wire [44:12] s12;
	wire [45:13] s13;
	wire [46:14] s14;
	wire [47:15] s15;
	wire [48:16] s16;
	wire [49:17] s17;
	wire [50:18] s18;
	wire [51:19] s19;
	wire [52:20] s20;
	wire [53:21] s21;
	wire [54:22] s22;
	wire [55:23] s23;
	wire [56:24] s24;
	wire [57:25] s25;
	wire [58:26] s26;
	wire [59:27] s27;
	wire [60:28] s28;
	wire [61:29] s29;
	wire [62:30] s30;
	wire [63:31] s31;

	assign s0[32] = zero;

	assign p0[31] = y[0]&x[31], p0[30] = y[0]&x[30], p0[29] = y[0]&x[29], p0[28] = y[0]&x[28], p0[27] = y[0]&x[27], p0[26] = y[0]&x[26], p0[25] = y[0]&x[25], p0[24] = y[0]&x[24], p0[23] = y[0]&x[23], p0[22] = y[0]&x[22], p0[21] = y[0]&x[21], p0[20] = y[0]&x[20], p0[19] = y[0]&x[19], p0[18] = y[0]&x[18], p0[17] = y[0]&x[17], p0[16] = y[0]&x[16], p0[15] = y[0]&x[15], p0[14] = y[0]&x[14], p0[13] = y[0]&x[13], p0[12] = y[0]&x[12], p0[11] = y[0]&x[11], p0[10] = y[0]&x[10], p0[9] = y[0]&x[9], p0[8] = y[0]&x[8], p0[7] = y[0]&x[7], p0[6] = y[0]&x[6], p0[5] = y[0]&x[5], p0[4] = y[0]&x[4], p0[3] = y[0]&x[3], p0[2] = y[0]&x[2], p0[1] = y[0]&x[1], p0[0] = y[0]&x[0];
	assign p1[32] = y[1]&x[31], p1[31] = y[1]&x[30], p1[30] = y[1]&x[29], p1[29] = y[1]&x[28], p1[28] = y[1]&x[27], p1[27] = y[1]&x[26], p1[26] = y[1]&x[25], p1[25] = y[1]&x[24], p1[24] = y[1]&x[23], p1[23] = y[1]&x[22], p1[22] = y[1]&x[21], p1[21] = y[1]&x[20], p1[20] = y[1]&x[19], p1[19] = y[1]&x[18], p1[18] = y[1]&x[17], p1[17] = y[1]&x[16], p1[16] = y[1]&x[15], p1[15] = y[1]&x[14], p1[14] = y[1]&x[13], p1[13] = y[1]&x[12], p1[12] = y[1]&x[11], p1[11] = y[1]&x[10], p1[10] = y[1]&x[9], p1[9] = y[1]&x[8], p1[8] = y[1]&x[7], p1[7] = y[1]&x[6], p1[6] = y[1]&x[5], p1[5] = y[1]&x[4], p1[4] = y[1]&x[3], p1[3] = y[1]&x[2], p1[2] = y[1]&x[1], p1[1] = y[1]&x[0];
	assign p2[33] = y[2]&x[31], p2[32] = y[2]&x[30], p2[31] = y[2]&x[29], p2[30] = y[2]&x[28], p2[29] = y[2]&x[27], p2[28] = y[2]&x[26], p2[27] = y[2]&x[25], p2[26] = y[2]&x[24], p2[25] = y[2]&x[23], p2[24] = y[2]&x[22], p2[23] = y[2]&x[21], p2[22] = y[2]&x[20], p2[21] = y[2]&x[19], p2[20] = y[2]&x[18], p2[19] = y[2]&x[17], p2[18] = y[2]&x[16], p2[17] = y[2]&x[15], p2[16] = y[2]&x[14], p2[15] = y[2]&x[13], p2[14] = y[2]&x[12], p2[13] = y[2]&x[11], p2[12] = y[2]&x[10], p2[11] = y[2]&x[9], p2[10] = y[2]&x[8], p2[9] = y[2]&x[7], p2[8] = y[2]&x[6], p2[7] = y[2]&x[5], p2[6] = y[2]&x[4], p2[5] = y[2]&x[3], p2[4] = y[2]&x[2], p2[3] = y[2]&x[1], p2[2] = y[2]&x[0];
	assign p3[34] = y[3]&x[31], p3[33] = y[3]&x[30], p3[32] = y[3]&x[29], p3[31] = y[3]&x[28], p3[30] = y[3]&x[27], p3[29] = y[3]&x[26], p3[28] = y[3]&x[25], p3[27] = y[3]&x[24], p3[26] = y[3]&x[23], p3[25] = y[3]&x[22], p3[24] = y[3]&x[21], p3[23] = y[3]&x[20], p3[22] = y[3]&x[19], p3[21] = y[3]&x[18], p3[20] = y[3]&x[17], p3[19] = y[3]&x[16], p3[18] = y[3]&x[15], p3[17] = y[3]&x[14], p3[16] = y[3]&x[13], p3[15] = y[3]&x[12], p3[14] = y[3]&x[11], p3[13] = y[3]&x[10], p3[12] = y[3]&x[9], p3[11] = y[3]&x[8], p3[10] = y[3]&x[7], p3[9] = y[3]&x[6], p3[8] = y[3]&x[5], p3[7] = y[3]&x[4], p3[6] = y[3]&x[3], p3[5] = y[3]&x[2], p3[4] = y[3]&x[1], p3[3] = y[3]&x[0];
	assign p4[35] = y[4]&x[31], p4[34] = y[4]&x[30], p4[33] = y[4]&x[29], p4[32] = y[4]&x[28], p4[31] = y[4]&x[27], p4[30] = y[4]&x[26], p4[29] = y[4]&x[25], p4[28] = y[4]&x[24], p4[27] = y[4]&x[23], p4[26] = y[4]&x[22], p4[25] = y[4]&x[21], p4[24] = y[4]&x[20], p4[23] = y[4]&x[19], p4[22] = y[4]&x[18], p4[21] = y[4]&x[17], p4[20] = y[4]&x[16], p4[19] = y[4]&x[15], p4[18] = y[4]&x[14], p4[17] = y[4]&x[13], p4[16] = y[4]&x[12], p4[15] = y[4]&x[11], p4[14] = y[4]&x[10], p4[13] = y[4]&x[9], p4[12] = y[4]&x[8], p4[11] = y[4]&x[7], p4[10] = y[4]&x[6], p4[9] = y[4]&x[5], p4[8] = y[4]&x[4], p4[7] = y[4]&x[3], p4[6] = y[4]&x[2], p4[5] = y[4]&x[1], p4[4] = y[4]&x[0];
	assign p5[36] = y[5]&x[31], p5[35] = y[5]&x[30], p5[34] = y[5]&x[29], p5[33] = y[5]&x[28], p5[32] = y[5]&x[27], p5[31] = y[5]&x[26], p5[30] = y[5]&x[25], p5[29] = y[5]&x[24], p5[28] = y[5]&x[23], p5[27] = y[5]&x[22], p5[26] = y[5]&x[21], p5[25] = y[5]&x[20], p5[24] = y[5]&x[19], p5[23] = y[5]&x[18], p5[22] = y[5]&x[17], p5[21] = y[5]&x[16], p5[20] = y[5]&x[15], p5[19] = y[5]&x[14], p5[18] = y[5]&x[13], p5[17] = y[5]&x[12], p5[16] = y[5]&x[11], p5[15] = y[5]&x[10], p5[14] = y[5]&x[9], p5[13] = y[5]&x[8], p5[12] = y[5]&x[7], p5[11] = y[5]&x[6], p5[10] = y[5]&x[5], p5[9] = y[5]&x[4], p5[8] = y[5]&x[3], p5[7] = y[5]&x[2], p5[6] = y[5]&x[1], p5[5] = y[5]&x[0];
	assign p6[37] = y[6]&x[31], p6[36] = y[6]&x[30], p6[35] = y[6]&x[29], p6[34] = y[6]&x[28], p6[33] = y[6]&x[27], p6[32] = y[6]&x[26], p6[31] = y[6]&x[25], p6[30] = y[6]&x[24], p6[29] = y[6]&x[23], p6[28] = y[6]&x[22], p6[27] = y[6]&x[21], p6[26] = y[6]&x[20], p6[25] = y[6]&x[19], p6[24] = y[6]&x[18], p6[23] = y[6]&x[17], p6[22] = y[6]&x[16], p6[21] = y[6]&x[15], p6[20] = y[6]&x[14], p6[19] = y[6]&x[13], p6[18] = y[6]&x[12], p6[17] = y[6]&x[11], p6[16] = y[6]&x[10], p6[15] = y[6]&x[9], p6[14] = y[6]&x[8], p6[13] = y[6]&x[7], p6[12] = y[6]&x[6], p6[11] = y[6]&x[5], p6[10] = y[6]&x[4], p6[9] = y[6]&x[3], p6[8] = y[6]&x[2], p6[7] = y[6]&x[1], p6[6] = y[6]&x[0];
	assign p7[38] = y[7]&x[31], p7[37] = y[7]&x[30], p7[36] = y[7]&x[29], p7[35] = y[7]&x[28], p7[34] = y[7]&x[27], p7[33] = y[7]&x[26], p7[32] = y[7]&x[25], p7[31] = y[7]&x[24], p7[30] = y[7]&x[23], p7[29] = y[7]&x[22], p7[28] = y[7]&x[21], p7[27] = y[7]&x[20], p7[26] = y[7]&x[19], p7[25] = y[7]&x[18], p7[24] = y[7]&x[17], p7[23] = y[7]&x[16], p7[22] = y[7]&x[15], p7[21] = y[7]&x[14], p7[20] = y[7]&x[13], p7[19] = y[7]&x[12], p7[18] = y[7]&x[11], p7[17] = y[7]&x[10], p7[16] = y[7]&x[9], p7[15] = y[7]&x[8], p7[14] = y[7]&x[7], p7[13] = y[7]&x[6], p7[12] = y[7]&x[5], p7[11] = y[7]&x[4], p7[10] = y[7]&x[3], p7[9] = y[7]&x[2], p7[8] = y[7]&x[1], p7[7] = y[7]&x[0];
	assign p8[39] = y[8]&x[31], p8[38] = y[8]&x[30], p8[37] = y[8]&x[29], p8[36] = y[8]&x[28], p8[35] = y[8]&x[27], p8[34] = y[8]&x[26], p8[33] = y[8]&x[25], p8[32] = y[8]&x[24], p8[31] = y[8]&x[23], p8[30] = y[8]&x[22], p8[29] = y[8]&x[21], p8[28] = y[8]&x[20], p8[27] = y[8]&x[19], p8[26] = y[8]&x[18], p8[25] = y[8]&x[17], p8[24] = y[8]&x[16], p8[23] = y[8]&x[15], p8[22] = y[8]&x[14], p8[21] = y[8]&x[13], p8[20] = y[8]&x[12], p8[19] = y[8]&x[11], p8[18] = y[8]&x[10], p8[17] = y[8]&x[9], p8[16] = y[8]&x[8], p8[15] = y[8]&x[7], p8[14] = y[8]&x[6], p8[13] = y[8]&x[5], p8[12] = y[8]&x[4], p8[11] = y[8]&x[3], p8[10] = y[8]&x[2], p8[9] = y[8]&x[1], p8[8] = y[8]&x[0];
	assign p9[40] = y[9]&x[31], p9[39] = y[9]&x[30], p9[38] = y[9]&x[29], p9[37] = y[9]&x[28], p9[36] = y[9]&x[27], p9[35] = y[9]&x[26], p9[34] = y[9]&x[25], p9[33] = y[9]&x[24], p9[32] = y[9]&x[23], p9[31] = y[9]&x[22], p9[30] = y[9]&x[21], p9[29] = y[9]&x[20], p9[28] = y[9]&x[19], p9[27] = y[9]&x[18], p9[26] = y[9]&x[17], p9[25] = y[9]&x[16], p9[24] = y[9]&x[15], p9[23] = y[9]&x[14], p9[22] = y[9]&x[13], p9[21] = y[9]&x[12], p9[20] = y[9]&x[11], p9[19] = y[9]&x[10], p9[18] = y[9]&x[9], p9[17] = y[9]&x[8], p9[16] = y[9]&x[7], p9[15] = y[9]&x[6], p9[14] = y[9]&x[5], p9[13] = y[9]&x[4], p9[12] = y[9]&x[3], p9[11] = y[9]&x[2], p9[10] = y[9]&x[1], p9[9] = y[9]&x[0];
	assign p10[41] = y[10]&x[31], p10[40] = y[10]&x[30], p10[39] = y[10]&x[29], p10[38] = y[10]&x[28], p10[37] = y[10]&x[27], p10[36] = y[10]&x[26], p10[35] = y[10]&x[25], p10[34] = y[10]&x[24], p10[33] = y[10]&x[23], p10[32] = y[10]&x[22], p10[31] = y[10]&x[21], p10[30] = y[10]&x[20], p10[29] = y[10]&x[19], p10[28] = y[10]&x[18], p10[27] = y[10]&x[17], p10[26] = y[10]&x[16], p10[25] = y[10]&x[15], p10[24] = y[10]&x[14], p10[23] = y[10]&x[13], p10[22] = y[10]&x[12], p10[21] = y[10]&x[11], p10[20] = y[10]&x[10], p10[19] = y[10]&x[9], p10[18] = y[10]&x[8], p10[17] = y[10]&x[7], p10[16] = y[10]&x[6], p10[15] = y[10]&x[5], p10[14] = y[10]&x[4], p10[13] = y[10]&x[3], p10[12] = y[10]&x[2], p10[11] = y[10]&x[1], p10[10] = y[10]&x[0];
	assign p11[42] = y[11]&x[31], p11[41] = y[11]&x[30], p11[40] = y[11]&x[29], p11[39] = y[11]&x[28], p11[38] = y[11]&x[27], p11[37] = y[11]&x[26], p11[36] = y[11]&x[25], p11[35] = y[11]&x[24], p11[34] = y[11]&x[23], p11[33] = y[11]&x[22], p11[32] = y[11]&x[21], p11[31] = y[11]&x[20], p11[30] = y[11]&x[19], p11[29] = y[11]&x[18], p11[28] = y[11]&x[17], p11[27] = y[11]&x[16], p11[26] = y[11]&x[15], p11[25] = y[11]&x[14], p11[24] = y[11]&x[13], p11[23] = y[11]&x[12], p11[22] = y[11]&x[11], p11[21] = y[11]&x[10], p11[20] = y[11]&x[9], p11[19] = y[11]&x[8], p11[18] = y[11]&x[7], p11[17] = y[11]&x[6], p11[16] = y[11]&x[5], p11[15] = y[11]&x[4], p11[14] = y[11]&x[3], p11[13] = y[11]&x[2], p11[12] = y[11]&x[1], p11[11] = y[11]&x[0];
	assign p12[43] = y[12]&x[31], p12[42] = y[12]&x[30], p12[41] = y[12]&x[29], p12[40] = y[12]&x[28], p12[39] = y[12]&x[27], p12[38] = y[12]&x[26], p12[37] = y[12]&x[25], p12[36] = y[12]&x[24], p12[35] = y[12]&x[23], p12[34] = y[12]&x[22], p12[33] = y[12]&x[21], p12[32] = y[12]&x[20], p12[31] = y[12]&x[19], p12[30] = y[12]&x[18], p12[29] = y[12]&x[17], p12[28] = y[12]&x[16], p12[27] = y[12]&x[15], p12[26] = y[12]&x[14], p12[25] = y[12]&x[13], p12[24] = y[12]&x[12], p12[23] = y[12]&x[11], p12[22] = y[12]&x[10], p12[21] = y[12]&x[9], p12[20] = y[12]&x[8], p12[19] = y[12]&x[7], p12[18] = y[12]&x[6], p12[17] = y[12]&x[5], p12[16] = y[12]&x[4], p12[15] = y[12]&x[3], p12[14] = y[12]&x[2], p12[13] = y[12]&x[1], p12[12] = y[12]&x[0];
	assign p13[44] = y[13]&x[31], p13[43] = y[13]&x[30], p13[42] = y[13]&x[29], p13[41] = y[13]&x[28], p13[40] = y[13]&x[27], p13[39] = y[13]&x[26], p13[38] = y[13]&x[25], p13[37] = y[13]&x[24], p13[36] = y[13]&x[23], p13[35] = y[13]&x[22], p13[34] = y[13]&x[21], p13[33] = y[13]&x[20], p13[32] = y[13]&x[19], p13[31] = y[13]&x[18], p13[30] = y[13]&x[17], p13[29] = y[13]&x[16], p13[28] = y[13]&x[15], p13[27] = y[13]&x[14], p13[26] = y[13]&x[13], p13[25] = y[13]&x[12], p13[24] = y[13]&x[11], p13[23] = y[13]&x[10], p13[22] = y[13]&x[9], p13[21] = y[13]&x[8], p13[20] = y[13]&x[7], p13[19] = y[13]&x[6], p13[18] = y[13]&x[5], p13[17] = y[13]&x[4], p13[16] = y[13]&x[3], p13[15] = y[13]&x[2], p13[14] = y[13]&x[1], p13[13] = y[13]&x[0];
	assign p14[45] = y[14]&x[31], p14[44] = y[14]&x[30], p14[43] = y[14]&x[29], p14[42] = y[14]&x[28], p14[41] = y[14]&x[27], p14[40] = y[14]&x[26], p14[39] = y[14]&x[25], p14[38] = y[14]&x[24], p14[37] = y[14]&x[23], p14[36] = y[14]&x[22], p14[35] = y[14]&x[21], p14[34] = y[14]&x[20], p14[33] = y[14]&x[19], p14[32] = y[14]&x[18], p14[31] = y[14]&x[17], p14[30] = y[14]&x[16], p14[29] = y[14]&x[15], p14[28] = y[14]&x[14], p14[27] = y[14]&x[13], p14[26] = y[14]&x[12], p14[25] = y[14]&x[11], p14[24] = y[14]&x[10], p14[23] = y[14]&x[9], p14[22] = y[14]&x[8], p14[21] = y[14]&x[7], p14[20] = y[14]&x[6], p14[19] = y[14]&x[5], p14[18] = y[14]&x[4], p14[17] = y[14]&x[3], p14[16] = y[14]&x[2], p14[15] = y[14]&x[1], p14[14] = y[14]&x[0];
	assign p15[46] = y[15]&x[31], p15[45] = y[15]&x[30], p15[44] = y[15]&x[29], p15[43] = y[15]&x[28], p15[42] = y[15]&x[27], p15[41] = y[15]&x[26], p15[40] = y[15]&x[25], p15[39] = y[15]&x[24], p15[38] = y[15]&x[23], p15[37] = y[15]&x[22], p15[36] = y[15]&x[21], p15[35] = y[15]&x[20], p15[34] = y[15]&x[19], p15[33] = y[15]&x[18], p15[32] = y[15]&x[17], p15[31] = y[15]&x[16], p15[30] = y[15]&x[15], p15[29] = y[15]&x[14], p15[28] = y[15]&x[13], p15[27] = y[15]&x[12], p15[26] = y[15]&x[11], p15[25] = y[15]&x[10], p15[24] = y[15]&x[9], p15[23] = y[15]&x[8], p15[22] = y[15]&x[7], p15[21] = y[15]&x[6], p15[20] = y[15]&x[5], p15[19] = y[15]&x[4], p15[18] = y[15]&x[3], p15[17] = y[15]&x[2], p15[16] = y[15]&x[1], p15[15] = y[15]&x[0];
	assign p16[47] = y[16]&x[31], p16[46] = y[16]&x[30], p16[45] = y[16]&x[29], p16[44] = y[16]&x[28], p16[43] = y[16]&x[27], p16[42] = y[16]&x[26], p16[41] = y[16]&x[25], p16[40] = y[16]&x[24], p16[39] = y[16]&x[23], p16[38] = y[16]&x[22], p16[37] = y[16]&x[21], p16[36] = y[16]&x[20], p16[35] = y[16]&x[19], p16[34] = y[16]&x[18], p16[33] = y[16]&x[17], p16[32] = y[16]&x[16], p16[31] = y[16]&x[15], p16[30] = y[16]&x[14], p16[29] = y[16]&x[13], p16[28] = y[16]&x[12], p16[27] = y[16]&x[11], p16[26] = y[16]&x[10], p16[25] = y[16]&x[9], p16[24] = y[16]&x[8], p16[23] = y[16]&x[7], p16[22] = y[16]&x[6], p16[21] = y[16]&x[5], p16[20] = y[16]&x[4], p16[19] = y[16]&x[3], p16[18] = y[16]&x[2], p16[17] = y[16]&x[1], p16[16] = y[16]&x[0];
	assign p17[48] = y[17]&x[31], p17[47] = y[17]&x[30], p17[46] = y[17]&x[29], p17[45] = y[17]&x[28], p17[44] = y[17]&x[27], p17[43] = y[17]&x[26], p17[42] = y[17]&x[25], p17[41] = y[17]&x[24], p17[40] = y[17]&x[23], p17[39] = y[17]&x[22], p17[38] = y[17]&x[21], p17[37] = y[17]&x[20], p17[36] = y[17]&x[19], p17[35] = y[17]&x[18], p17[34] = y[17]&x[17], p17[33] = y[17]&x[16], p17[32] = y[17]&x[15], p17[31] = y[17]&x[14], p17[30] = y[17]&x[13], p17[29] = y[17]&x[12], p17[28] = y[17]&x[11], p17[27] = y[17]&x[10], p17[26] = y[17]&x[9], p17[25] = y[17]&x[8], p17[24] = y[17]&x[7], p17[23] = y[17]&x[6], p17[22] = y[17]&x[5], p17[21] = y[17]&x[4], p17[20] = y[17]&x[3], p17[19] = y[17]&x[2], p17[18] = y[17]&x[1], p17[17] = y[17]&x[0];
	assign p18[49] = y[18]&x[31], p18[48] = y[18]&x[30], p18[47] = y[18]&x[29], p18[46] = y[18]&x[28], p18[45] = y[18]&x[27], p18[44] = y[18]&x[26], p18[43] = y[18]&x[25], p18[42] = y[18]&x[24], p18[41] = y[18]&x[23], p18[40] = y[18]&x[22], p18[39] = y[18]&x[21], p18[38] = y[18]&x[20], p18[37] = y[18]&x[19], p18[36] = y[18]&x[18], p18[35] = y[18]&x[17], p18[34] = y[18]&x[16], p18[33] = y[18]&x[15], p18[32] = y[18]&x[14], p18[31] = y[18]&x[13], p18[30] = y[18]&x[12], p18[29] = y[18]&x[11], p18[28] = y[18]&x[10], p18[27] = y[18]&x[9], p18[26] = y[18]&x[8], p18[25] = y[18]&x[7], p18[24] = y[18]&x[6], p18[23] = y[18]&x[5], p18[22] = y[18]&x[4], p18[21] = y[18]&x[3], p18[20] = y[18]&x[2], p18[19] = y[18]&x[1], p18[18] = y[18]&x[0];
	assign p19[50] = y[19]&x[31], p19[49] = y[19]&x[30], p19[48] = y[19]&x[29], p19[47] = y[19]&x[28], p19[46] = y[19]&x[27], p19[45] = y[19]&x[26], p19[44] = y[19]&x[25], p19[43] = y[19]&x[24], p19[42] = y[19]&x[23], p19[41] = y[19]&x[22], p19[40] = y[19]&x[21], p19[39] = y[19]&x[20], p19[38] = y[19]&x[19], p19[37] = y[19]&x[18], p19[36] = y[19]&x[17], p19[35] = y[19]&x[16], p19[34] = y[19]&x[15], p19[33] = y[19]&x[14], p19[32] = y[19]&x[13], p19[31] = y[19]&x[12], p19[30] = y[19]&x[11], p19[29] = y[19]&x[10], p19[28] = y[19]&x[9], p19[27] = y[19]&x[8], p19[26] = y[19]&x[7], p19[25] = y[19]&x[6], p19[24] = y[19]&x[5], p19[23] = y[19]&x[4], p19[22] = y[19]&x[3], p19[21] = y[19]&x[2], p19[20] = y[19]&x[1], p19[19] = y[19]&x[0];
	assign p20[51] = y[20]&x[31], p20[50] = y[20]&x[30], p20[49] = y[20]&x[29], p20[48] = y[20]&x[28], p20[47] = y[20]&x[27], p20[46] = y[20]&x[26], p20[45] = y[20]&x[25], p20[44] = y[20]&x[24], p20[43] = y[20]&x[23], p20[42] = y[20]&x[22], p20[41] = y[20]&x[21], p20[40] = y[20]&x[20], p20[39] = y[20]&x[19], p20[38] = y[20]&x[18], p20[37] = y[20]&x[17], p20[36] = y[20]&x[16], p20[35] = y[20]&x[15], p20[34] = y[20]&x[14], p20[33] = y[20]&x[13], p20[32] = y[20]&x[12], p20[31] = y[20]&x[11], p20[30] = y[20]&x[10], p20[29] = y[20]&x[9], p20[28] = y[20]&x[8], p20[27] = y[20]&x[7], p20[26] = y[20]&x[6], p20[25] = y[20]&x[5], p20[24] = y[20]&x[4], p20[23] = y[20]&x[3], p20[22] = y[20]&x[2], p20[21] = y[20]&x[1], p20[20] = y[20]&x[0];
	assign p21[52] = y[21]&x[31], p21[51] = y[21]&x[30], p21[50] = y[21]&x[29], p21[49] = y[21]&x[28], p21[48] = y[21]&x[27], p21[47] = y[21]&x[26], p21[46] = y[21]&x[25], p21[45] = y[21]&x[24], p21[44] = y[21]&x[23], p21[43] = y[21]&x[22], p21[42] = y[21]&x[21], p21[41] = y[21]&x[20], p21[40] = y[21]&x[19], p21[39] = y[21]&x[18], p21[38] = y[21]&x[17], p21[37] = y[21]&x[16], p21[36] = y[21]&x[15], p21[35] = y[21]&x[14], p21[34] = y[21]&x[13], p21[33] = y[21]&x[12], p21[32] = y[21]&x[11], p21[31] = y[21]&x[10], p21[30] = y[21]&x[9], p21[29] = y[21]&x[8], p21[28] = y[21]&x[7], p21[27] = y[21]&x[6], p21[26] = y[21]&x[5], p21[25] = y[21]&x[4], p21[24] = y[21]&x[3], p21[23] = y[21]&x[2], p21[22] = y[21]&x[1], p21[21] = y[21]&x[0];
	assign p22[53] = y[22]&x[31], p22[52] = y[22]&x[30], p22[51] = y[22]&x[29], p22[50] = y[22]&x[28], p22[49] = y[22]&x[27], p22[48] = y[22]&x[26], p22[47] = y[22]&x[25], p22[46] = y[22]&x[24], p22[45] = y[22]&x[23], p22[44] = y[22]&x[22], p22[43] = y[22]&x[21], p22[42] = y[22]&x[20], p22[41] = y[22]&x[19], p22[40] = y[22]&x[18], p22[39] = y[22]&x[17], p22[38] = y[22]&x[16], p22[37] = y[22]&x[15], p22[36] = y[22]&x[14], p22[35] = y[22]&x[13], p22[34] = y[22]&x[12], p22[33] = y[22]&x[11], p22[32] = y[22]&x[10], p22[31] = y[22]&x[9], p22[30] = y[22]&x[8], p22[29] = y[22]&x[7], p22[28] = y[22]&x[6], p22[27] = y[22]&x[5], p22[26] = y[22]&x[4], p22[25] = y[22]&x[3], p22[24] = y[22]&x[2], p22[23] = y[22]&x[1], p22[22] = y[22]&x[0];
	assign p23[54] = y[23]&x[31], p23[53] = y[23]&x[30], p23[52] = y[23]&x[29], p23[51] = y[23]&x[28], p23[50] = y[23]&x[27], p23[49] = y[23]&x[26], p23[48] = y[23]&x[25], p23[47] = y[23]&x[24], p23[46] = y[23]&x[23], p23[45] = y[23]&x[22], p23[44] = y[23]&x[21], p23[43] = y[23]&x[20], p23[42] = y[23]&x[19], p23[41] = y[23]&x[18], p23[40] = y[23]&x[17], p23[39] = y[23]&x[16], p23[38] = y[23]&x[15], p23[37] = y[23]&x[14], p23[36] = y[23]&x[13], p23[35] = y[23]&x[12], p23[34] = y[23]&x[11], p23[33] = y[23]&x[10], p23[32] = y[23]&x[9], p23[31] = y[23]&x[8], p23[30] = y[23]&x[7], p23[29] = y[23]&x[6], p23[28] = y[23]&x[5], p23[27] = y[23]&x[4], p23[26] = y[23]&x[3], p23[25] = y[23]&x[2], p23[24] = y[23]&x[1], p23[23] = y[23]&x[0];
	assign p24[55] = y[24]&x[31], p24[54] = y[24]&x[30], p24[53] = y[24]&x[29], p24[52] = y[24]&x[28], p24[51] = y[24]&x[27], p24[50] = y[24]&x[26], p24[49] = y[24]&x[25], p24[48] = y[24]&x[24], p24[47] = y[24]&x[23], p24[46] = y[24]&x[22], p24[45] = y[24]&x[21], p24[44] = y[24]&x[20], p24[43] = y[24]&x[19], p24[42] = y[24]&x[18], p24[41] = y[24]&x[17], p24[40] = y[24]&x[16], p24[39] = y[24]&x[15], p24[38] = y[24]&x[14], p24[37] = y[24]&x[13], p24[36] = y[24]&x[12], p24[35] = y[24]&x[11], p24[34] = y[24]&x[10], p24[33] = y[24]&x[9], p24[32] = y[24]&x[8], p24[31] = y[24]&x[7], p24[30] = y[24]&x[6], p24[29] = y[24]&x[5], p24[28] = y[24]&x[4], p24[27] = y[24]&x[3], p24[26] = y[24]&x[2], p24[25] = y[24]&x[1], p24[24] = y[24]&x[0];
	assign p25[56] = y[25]&x[31], p25[55] = y[25]&x[30], p25[54] = y[25]&x[29], p25[53] = y[25]&x[28], p25[52] = y[25]&x[27], p25[51] = y[25]&x[26], p25[50] = y[25]&x[25], p25[49] = y[25]&x[24], p25[48] = y[25]&x[23], p25[47] = y[25]&x[22], p25[46] = y[25]&x[21], p25[45] = y[25]&x[20], p25[44] = y[25]&x[19], p25[43] = y[25]&x[18], p25[42] = y[25]&x[17], p25[41] = y[25]&x[16], p25[40] = y[25]&x[15], p25[39] = y[25]&x[14], p25[38] = y[25]&x[13], p25[37] = y[25]&x[12], p25[36] = y[25]&x[11], p25[35] = y[25]&x[10], p25[34] = y[25]&x[9], p25[33] = y[25]&x[8], p25[32] = y[25]&x[7], p25[31] = y[25]&x[6], p25[30] = y[25]&x[5], p25[29] = y[25]&x[4], p25[28] = y[25]&x[3], p25[27] = y[25]&x[2], p25[26] = y[25]&x[1], p25[25] = y[25]&x[0];
	assign p26[57] = y[26]&x[31], p26[56] = y[26]&x[30], p26[55] = y[26]&x[29], p26[54] = y[26]&x[28], p26[53] = y[26]&x[27], p26[52] = y[26]&x[26], p26[51] = y[26]&x[25], p26[50] = y[26]&x[24], p26[49] = y[26]&x[23], p26[48] = y[26]&x[22], p26[47] = y[26]&x[21], p26[46] = y[26]&x[20], p26[45] = y[26]&x[19], p26[44] = y[26]&x[18], p26[43] = y[26]&x[17], p26[42] = y[26]&x[16], p26[41] = y[26]&x[15], p26[40] = y[26]&x[14], p26[39] = y[26]&x[13], p26[38] = y[26]&x[12], p26[37] = y[26]&x[11], p26[36] = y[26]&x[10], p26[35] = y[26]&x[9], p26[34] = y[26]&x[8], p26[33] = y[26]&x[7], p26[32] = y[26]&x[6], p26[31] = y[26]&x[5], p26[30] = y[26]&x[4], p26[29] = y[26]&x[3], p26[28] = y[26]&x[2], p26[27] = y[26]&x[1], p26[26] = y[26]&x[0];
	assign p27[58] = y[27]&x[31], p27[57] = y[27]&x[30], p27[56] = y[27]&x[29], p27[55] = y[27]&x[28], p27[54] = y[27]&x[27], p27[53] = y[27]&x[26], p27[52] = y[27]&x[25], p27[51] = y[27]&x[24], p27[50] = y[27]&x[23], p27[49] = y[27]&x[22], p27[48] = y[27]&x[21], p27[47] = y[27]&x[20], p27[46] = y[27]&x[19], p27[45] = y[27]&x[18], p27[44] = y[27]&x[17], p27[43] = y[27]&x[16], p27[42] = y[27]&x[15], p27[41] = y[27]&x[14], p27[40] = y[27]&x[13], p27[39] = y[27]&x[12], p27[38] = y[27]&x[11], p27[37] = y[27]&x[10], p27[36] = y[27]&x[9], p27[35] = y[27]&x[8], p27[34] = y[27]&x[7], p27[33] = y[27]&x[6], p27[32] = y[27]&x[5], p27[31] = y[27]&x[4], p27[30] = y[27]&x[3], p27[29] = y[27]&x[2], p27[28] = y[27]&x[1], p27[27] = y[27]&x[0];
	assign p28[59] = y[28]&x[31], p28[58] = y[28]&x[30], p28[57] = y[28]&x[29], p28[56] = y[28]&x[28], p28[55] = y[28]&x[27], p28[54] = y[28]&x[26], p28[53] = y[28]&x[25], p28[52] = y[28]&x[24], p28[51] = y[28]&x[23], p28[50] = y[28]&x[22], p28[49] = y[28]&x[21], p28[48] = y[28]&x[20], p28[47] = y[28]&x[19], p28[46] = y[28]&x[18], p28[45] = y[28]&x[17], p28[44] = y[28]&x[16], p28[43] = y[28]&x[15], p28[42] = y[28]&x[14], p28[41] = y[28]&x[13], p28[40] = y[28]&x[12], p28[39] = y[28]&x[11], p28[38] = y[28]&x[10], p28[37] = y[28]&x[9], p28[36] = y[28]&x[8], p28[35] = y[28]&x[7], p28[34] = y[28]&x[6], p28[33] = y[28]&x[5], p28[32] = y[28]&x[4], p28[31] = y[28]&x[3], p28[30] = y[28]&x[2], p28[29] = y[28]&x[1], p28[28] = y[28]&x[0];
	assign p29[60] = y[29]&x[31], p29[59] = y[29]&x[30], p29[58] = y[29]&x[29], p29[57] = y[29]&x[28], p29[56] = y[29]&x[27], p29[55] = y[29]&x[26], p29[54] = y[29]&x[25], p29[53] = y[29]&x[24], p29[52] = y[29]&x[23], p29[51] = y[29]&x[22], p29[50] = y[29]&x[21], p29[49] = y[29]&x[20], p29[48] = y[29]&x[19], p29[47] = y[29]&x[18], p29[46] = y[29]&x[17], p29[45] = y[29]&x[16], p29[44] = y[29]&x[15], p29[43] = y[29]&x[14], p29[42] = y[29]&x[13], p29[41] = y[29]&x[12], p29[40] = y[29]&x[11], p29[39] = y[29]&x[10], p29[38] = y[29]&x[9], p29[37] = y[29]&x[8], p29[36] = y[29]&x[7], p29[35] = y[29]&x[6], p29[34] = y[29]&x[5], p29[33] = y[29]&x[4], p29[32] = y[29]&x[3], p29[31] = y[29]&x[2], p29[30] = y[29]&x[1], p29[29] = y[29]&x[0];
	assign p30[61] = y[30]&x[31], p30[60] = y[30]&x[30], p30[59] = y[30]&x[29], p30[58] = y[30]&x[28], p30[57] = y[30]&x[27], p30[56] = y[30]&x[26], p30[55] = y[30]&x[25], p30[54] = y[30]&x[24], p30[53] = y[30]&x[23], p30[52] = y[30]&x[22], p30[51] = y[30]&x[21], p30[50] = y[30]&x[20], p30[49] = y[30]&x[19], p30[48] = y[30]&x[18], p30[47] = y[30]&x[17], p30[46] = y[30]&x[16], p30[45] = y[30]&x[15], p30[44] = y[30]&x[14], p30[43] = y[30]&x[13], p30[42] = y[30]&x[12], p30[41] = y[30]&x[11], p30[40] = y[30]&x[10], p30[39] = y[30]&x[9], p30[38] = y[30]&x[8], p30[37] = y[30]&x[7], p30[36] = y[30]&x[6], p30[35] = y[30]&x[5], p30[34] = y[30]&x[4], p30[33] = y[30]&x[3], p30[32] = y[30]&x[2], p30[31] = y[30]&x[1], p30[30] = y[30]&x[0];
	assign p31[62] = y[31]&x[31], p31[61] = y[31]&x[30], p31[60] = y[31]&x[29], p31[59] = y[31]&x[28], p31[58] = y[31]&x[27], p31[57] = y[31]&x[26], p31[56] = y[31]&x[25], p31[55] = y[31]&x[24], p31[54] = y[31]&x[23], p31[53] = y[31]&x[22], p31[52] = y[31]&x[21], p31[51] = y[31]&x[20], p31[50] = y[31]&x[19], p31[49] = y[31]&x[18], p31[48] = y[31]&x[17], p31[47] = y[31]&x[16], p31[46] = y[31]&x[15], p31[45] = y[31]&x[14], p31[44] = y[31]&x[13], p31[43] = y[31]&x[12], p31[42] = y[31]&x[11], p31[41] = y[31]&x[10], p31[40] = y[31]&x[9], p31[39] = y[31]&x[8], p31[38] = y[31]&x[7], p31[37] = y[31]&x[6], p31[36] = y[31]&x[5], p31[35] = y[31]&x[4], p31[34] = y[31]&x[3], p31[33] = y[31]&x[2], p31[32] = y[31]&x[1], p31[31] = y[31]&x[0];


	assign s0[31:0] = p0;

	Prefix_Add32 f1(s0[32:1], p1[32:1], zero, s1[32:1], s1[33]);
	Prefix_Add32 f2(s1[33:2], p2[33:2], zero, s2[33:2], s2[34]);
	Prefix_Add32 f3(s2[34:3], p3[34:3], zero, s3[34:3], s3[35]);
	Prefix_Add32 f4(s3[35:4], p4[35:4], zero, s4[35:4], s4[36]);
	Prefix_Add32 f5(s4[36:5], p5[36:5], zero, s5[36:5], s5[37]);
	Prefix_Add32 f6(s5[37:6], p6[37:6], zero, s6[37:6], s6[38]);
	Prefix_Add32 f7(s6[38:7], p7[38:7], zero, s7[38:7], s7[39]);
	Prefix_Add32 f8(s7[39:8], p8[39:8], zero, s8[39:8], s8[40]);
	Prefix_Add32 f9(s8[40:9], p9[40:9], zero, s9[40:9], s9[41]);
	Prefix_Add32 f10(s9[41:10], p10[41:10], zero, s10[41:10], s10[42]);
	Prefix_Add32 f11(s10[42:11], p11[42:11], zero, s11[42:11], s11[43]);
	Prefix_Add32 f12(s11[43:12], p12[43:12], zero, s12[43:12], s12[44]);
	Prefix_Add32 f13(s12[44:13], p13[44:13], zero, s13[44:13], s13[45]);
	Prefix_Add32 f14(s13[45:14], p14[45:14], zero, s14[45:14], s14[46]);
	Prefix_Add32 f15(s14[46:15], p15[46:15], zero, s15[46:15], s15[47]);
	Prefix_Add32 f16(s15[47:16], p16[47:16], zero, s16[47:16], s16[48]);
	Prefix_Add32 f17(s16[48:17], p17[48:17], zero, s17[48:17], s17[49]);
	Prefix_Add32 f18(s17[49:18], p18[49:18], zero, s18[49:18], s18[50]);
	Prefix_Add32 f19(s18[50:19], p19[50:19], zero, s19[50:19], s19[51]);
	Prefix_Add32 f20(s19[51:20], p20[51:20], zero, s20[51:20], s20[52]);
	Prefix_Add32 f21(s20[52:21], p21[52:21], zero, s21[52:21], s21[53]);
	Prefix_Add32 f22(s21[53:22], p22[53:22], zero, s22[53:22], s22[54]);
	Prefix_Add32 f23(s22[54:23], p23[54:23], zero, s23[54:23], s23[55]);
	Prefix_Add32 f24(s23[55:24], p24[55:24], zero, s24[55:24], s24[56]);
	Prefix_Add32 f25(s24[56:25], p25[56:25], zero, s25[56:25], s25[57]);
	Prefix_Add32 f26(s25[57:26], p26[57:26], zero, s26[57:26], s26[58]);
	Prefix_Add32 f27(s26[58:27], p27[58:27], zero, s27[58:27], s27[59]);
	Prefix_Add32 f28(s27[59:28], p28[59:28], zero, s28[59:28], s28[60]);
	Prefix_Add32 f29(s28[60:29], p29[60:29], zero, s29[60:29], s29[61]);
	Prefix_Add32 f30(s29[61:30], p30[61:30], zero, s30[61:30], s30[62]);
	Prefix_Add32 f31(s30[62:31], p31[62:31], zero, s31[62:31], s31[63]);


	assign P[0] = s0[0];
	assign P[1] = s1[1];
	assign P[2] = s2[2];
	assign P[3] = s3[3];
	assign P[4] = s4[4];
	assign P[5] = s5[5];
	assign P[6] = s6[6];
	assign P[7] = s7[7];
	assign P[8] = s8[8];
	assign P[9] = s9[9];
	assign P[10] = s10[10];
	assign P[11] = s11[11];
	assign P[12] = s12[12];
	assign P[13] = s13[13];
	assign P[14] = s14[14];
	assign P[15] = s15[15];
	assign P[16] = s16[16];
	assign P[17] = s17[17];
	assign P[18] = s18[18];
	assign P[19] = s19[19];
	assign P[20] = s20[20];
	assign P[21] = s21[21];
	assign P[22] = s22[22];
	assign P[23] = s23[23];
	assign P[24] = s24[24];
	assign P[25] = s25[25];
	assign P[26] = s26[26];
	assign P[27] = s27[27];
	assign P[28] = s28[28];
	assign P[29] = s29[29];
	assign P[30] = s30[30];

	assign P[63:31] = s31[63:31];


endmodule
