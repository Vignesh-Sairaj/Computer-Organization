module Prefix_Add32(x, y, cIn, s, cOut);

	input [31:0] x, y;
	input cIn;

	output [31:0] s;
	output cOut;

	wire [31:0] g0, p0, g1, p1, g2, p2, g3, p3, g4, p4, g5, p5;
	wire [32:0] c;

	assign g0[31:1] = x[31:1]&y[31:1];
	assign p0[31:0] = x^y;
	assign c[0] = cIn;
	assign g0[0] = x[0]&y[0] | c[0]&(x[0] | y[0]);



	assign g1[31] = g0[31] | p0[31]&g0[30], g1[30] = g0[30] | p0[30]&g0[29], g1[29] = g0[29] | p0[29]&g0[28], g1[28] = g0[28] | p0[28]&g0[27], g1[27] = g0[27] | p0[27]&g0[26], g1[26] = g0[26] | p0[26]&g0[25], g1[25] = g0[25] | p0[25]&g0[24], g1[24] = g0[24] | p0[24]&g0[23], g1[23] = g0[23] | p0[23]&g0[22], g1[22] = g0[22] | p0[22]&g0[21], g1[21] = g0[21] | p0[21]&g0[20], g1[20] = g0[20] | p0[20]&g0[19], g1[19] = g0[19] | p0[19]&g0[18], g1[18] = g0[18] | p0[18]&g0[17], g1[17] = g0[17] | p0[17]&g0[16], g1[16] = g0[16] | p0[16]&g0[15], g1[15] = g0[15] | p0[15]&g0[14], g1[14] = g0[14] | p0[14]&g0[13], g1[13] = g0[13] | p0[13]&g0[12], g1[12] = g0[12] | p0[12]&g0[11], g1[11] = g0[11] | p0[11]&g0[10], g1[10] = g0[10] | p0[10]&g0[9], g1[9] = g0[9] | p0[9]&g0[8], g1[8] = g0[8] | p0[8]&g0[7], g1[7] = g0[7] | p0[7]&g0[6], g1[6] = g0[6] | p0[6]&g0[5], g1[5] = g0[5] | p0[5]&g0[4], g1[4] = g0[4] | p0[4]&g0[3], g1[3] = g0[3] | p0[3]&g0[2], g1[2] = g0[2] | p0[2]&g0[1], g1[1] = g0[1] | p0[1]&g0[0], g1[0] = g0[0];
	assign p1[31] = p0[31]&p0[30], p1[30] = p0[30]&p0[29], p1[29] = p0[29]&p0[28], p1[28] = p0[28]&p0[27], p1[27] = p0[27]&p0[26], p1[26] = p0[26]&p0[25], p1[25] = p0[25]&p0[24], p1[24] = p0[24]&p0[23], p1[23] = p0[23]&p0[22], p1[22] = p0[22]&p0[21], p1[21] = p0[21]&p0[20], p1[20] = p0[20]&p0[19], p1[19] = p0[19]&p0[18], p1[18] = p0[18]&p0[17], p1[17] = p0[17]&p0[16], p1[16] = p0[16]&p0[15], p1[15] = p0[15]&p0[14], p1[14] = p0[14]&p0[13], p1[13] = p0[13]&p0[12], p1[12] = p0[12]&p0[11], p1[11] = p0[11]&p0[10], p1[10] = p0[10]&p0[9], p1[9] = p0[9]&p0[8], p1[8] = p0[8]&p0[7], p1[7] = p0[7]&p0[6], p1[6] = p0[6]&p0[5], p1[5] = p0[5]&p0[4], p1[4] = p0[4]&p0[3], p1[3] = p0[3]&p0[2], p1[2] = p0[2]&p0[1], p1[1] = p0[1]&p0[0], p1[0] = p0[0];

	assign g2[31] = g1[31] | p1[31]&g1[29], g2[30] = g1[30] | p1[30]&g1[28], g2[29] = g1[29] | p1[29]&g1[27], g2[28] = g1[28] | p1[28]&g1[26], g2[27] = g1[27] | p1[27]&g1[25], g2[26] = g1[26] | p1[26]&g1[24], g2[25] = g1[25] | p1[25]&g1[23], g2[24] = g1[24] | p1[24]&g1[22], g2[23] = g1[23] | p1[23]&g1[21], g2[22] = g1[22] | p1[22]&g1[20], g2[21] = g1[21] | p1[21]&g1[19], g2[20] = g1[20] | p1[20]&g1[18], g2[19] = g1[19] | p1[19]&g1[17], g2[18] = g1[18] | p1[18]&g1[16], g2[17] = g1[17] | p1[17]&g1[15], g2[16] = g1[16] | p1[16]&g1[14], g2[15] = g1[15] | p1[15]&g1[13], g2[14] = g1[14] | p1[14]&g1[12], g2[13] = g1[13] | p1[13]&g1[11], g2[12] = g1[12] | p1[12]&g1[10], g2[11] = g1[11] | p1[11]&g1[9], g2[10] = g1[10] | p1[10]&g1[8], g2[9] = g1[9] | p1[9]&g1[7], g2[8] = g1[8] | p1[8]&g1[6], g2[7] = g1[7] | p1[7]&g1[5], g2[6] = g1[6] | p1[6]&g1[4], g2[5] = g1[5] | p1[5]&g1[3], g2[4] = g1[4] | p1[4]&g1[2], g2[3] = g1[3] | p1[3]&g1[1], g2[2] = g1[2] | p1[2]&g1[0], g2[1] = g1[1], g2[0] = g1[0];
	assign p2[31] = p1[31]&p1[29], p2[30] = p1[30]&p1[28], p2[29] = p1[29]&p1[27], p2[28] = p1[28]&p1[26], p2[27] = p1[27]&p1[25], p2[26] = p1[26]&p1[24], p2[25] = p1[25]&p1[23], p2[24] = p1[24]&p1[22], p2[23] = p1[23]&p1[21], p2[22] = p1[22]&p1[20], p2[21] = p1[21]&p1[19], p2[20] = p1[20]&p1[18], p2[19] = p1[19]&p1[17], p2[18] = p1[18]&p1[16], p2[17] = p1[17]&p1[15], p2[16] = p1[16]&p1[14], p2[15] = p1[15]&p1[13], p2[14] = p1[14]&p1[12], p2[13] = p1[13]&p1[11], p2[12] = p1[12]&p1[10], p2[11] = p1[11]&p1[9], p2[10] = p1[10]&p1[8], p2[9] = p1[9]&p1[7], p2[8] = p1[8]&p1[6], p2[7] = p1[7]&p1[5], p2[6] = p1[6]&p1[4], p2[5] = p1[5]&p1[3], p2[4] = p1[4]&p1[2], p2[3] = p1[3]&p1[1], p2[2] = p1[2]&p1[0], p2[1] = p1[1], p2[0] = p1[0];

	assign g3[31] = g2[31] | p2[31]&g2[27], g3[30] = g2[30] | p2[30]&g2[26], g3[29] = g2[29] | p2[29]&g2[25], g3[28] = g2[28] | p2[28]&g2[24], g3[27] = g2[27] | p2[27]&g2[23], g3[26] = g2[26] | p2[26]&g2[22], g3[25] = g2[25] | p2[25]&g2[21], g3[24] = g2[24] | p2[24]&g2[20], g3[23] = g2[23] | p2[23]&g2[19], g3[22] = g2[22] | p2[22]&g2[18], g3[21] = g2[21] | p2[21]&g2[17], g3[20] = g2[20] | p2[20]&g2[16], g3[19] = g2[19] | p2[19]&g2[15], g3[18] = g2[18] | p2[18]&g2[14], g3[17] = g2[17] | p2[17]&g2[13], g3[16] = g2[16] | p2[16]&g2[12], g3[15] = g2[15] | p2[15]&g2[11], g3[14] = g2[14] | p2[14]&g2[10], g3[13] = g2[13] | p2[13]&g2[9], g3[12] = g2[12] | p2[12]&g2[8], g3[11] = g2[11] | p2[11]&g2[7], g3[10] = g2[10] | p2[10]&g2[6], g3[9] = g2[9] | p2[9]&g2[5], g3[8] = g2[8] | p2[8]&g2[4], g3[7] = g2[7] | p2[7]&g2[3], g3[6] = g2[6] | p2[6]&g2[2], g3[5] = g2[5] | p2[5]&g2[1], g3[4] = g2[4] | p2[4]&g2[0], g3[3] = g2[3], g3[2] = g2[2], g3[1] = g2[1], g3[0] = g2[0];
	assign p3[31] = p2[31]&p2[27], p3[30] = p2[30]&p2[26], p3[29] = p2[29]&p2[25], p3[28] = p2[28]&p2[24], p3[27] = p2[27]&p2[23], p3[26] = p2[26]&p2[22], p3[25] = p2[25]&p2[21], p3[24] = p2[24]&p2[20], p3[23] = p2[23]&p2[19], p3[22] = p2[22]&p2[18], p3[21] = p2[21]&p2[17], p3[20] = p2[20]&p2[16], p3[19] = p2[19]&p2[15], p3[18] = p2[18]&p2[14], p3[17] = p2[17]&p2[13], p3[16] = p2[16]&p2[12], p3[15] = p2[15]&p2[11], p3[14] = p2[14]&p2[10], p3[13] = p2[13]&p2[9], p3[12] = p2[12]&p2[8], p3[11] = p2[11]&p2[7], p3[10] = p2[10]&p2[6], p3[9] = p2[9]&p2[5], p3[8] = p2[8]&p2[4], p3[7] = p2[7]&p2[3], p3[6] = p2[6]&p2[2], p3[5] = p2[5]&p2[1], p3[4] = p2[4]&p2[0], p3[3] = p2[3], p3[2] = p2[2], p3[1] = p2[1], p3[0] = p2[0];

	assign g4[31] = g3[31] | p3[31]&g3[23], g4[30] = g3[30] | p3[30]&g3[22], g4[29] = g3[29] | p3[29]&g3[21], g4[28] = g3[28] | p3[28]&g3[20], g4[27] = g3[27] | p3[27]&g3[19], g4[26] = g3[26] | p3[26]&g3[18], g4[25] = g3[25] | p3[25]&g3[17], g4[24] = g3[24] | p3[24]&g3[16], g4[23] = g3[23] | p3[23]&g3[15], g4[22] = g3[22] | p3[22]&g3[14], g4[21] = g3[21] | p3[21]&g3[13], g4[20] = g3[20] | p3[20]&g3[12], g4[19] = g3[19] | p3[19]&g3[11], g4[18] = g3[18] | p3[18]&g3[10], g4[17] = g3[17] | p3[17]&g3[9], g4[16] = g3[16] | p3[16]&g3[8], g4[15] = g3[15] | p3[15]&g3[7], g4[14] = g3[14] | p3[14]&g3[6], g4[13] = g3[13] | p3[13]&g3[5], g4[12] = g3[12] | p3[12]&g3[4], g4[11] = g3[11] | p3[11]&g3[3], g4[10] = g3[10] | p3[10]&g3[2], g4[9] = g3[9] | p3[9]&g3[1], g4[8] = g3[8] | p3[8]&g3[0], g4[7] = g3[7], g4[6] = g3[6], g4[5] = g3[5], g4[4] = g3[4], g4[3] = g3[3], g4[2] = g3[2], g4[1] = g3[1], g4[0] = g3[0];
	assign p4[31] = p3[31]&p3[23], p4[30] = p3[30]&p3[22], p4[29] = p3[29]&p3[21], p4[28] = p3[28]&p3[20], p4[27] = p3[27]&p3[19], p4[26] = p3[26]&p3[18], p4[25] = p3[25]&p3[17], p4[24] = p3[24]&p3[16], p4[23] = p3[23]&p3[15], p4[22] = p3[22]&p3[14], p4[21] = p3[21]&p3[13], p4[20] = p3[20]&p3[12], p4[19] = p3[19]&p3[11], p4[18] = p3[18]&p3[10], p4[17] = p3[17]&p3[9], p4[16] = p3[16]&p3[8], p4[15] = p3[15]&p3[7], p4[14] = p3[14]&p3[6], p4[13] = p3[13]&p3[5], p4[12] = p3[12]&p3[4], p4[11] = p3[11]&p3[3], p4[10] = p3[10]&p3[2], p4[9] = p3[9]&p3[1], p4[8] = p3[8]&p3[0], p4[7] = p3[7], p4[6] = p3[6], p4[5] = p3[5], p4[4] = p3[4], p4[3] = p3[3], p4[2] = p3[2], p4[1] = p3[1], p4[0] = p3[0];

	assign g5[31] = g4[31] | p4[31]&g4[15], g5[30] = g4[30] | p4[30]&g4[14], g5[29] = g4[29] | p4[29]&g4[13], g5[28] = g4[28] | p4[28]&g4[12], g5[27] = g4[27] | p4[27]&g4[11], g5[26] = g4[26] | p4[26]&g4[10], g5[25] = g4[25] | p4[25]&g4[9], g5[24] = g4[24] | p4[24]&g4[8], g5[23] = g4[23] | p4[23]&g4[7], g5[22] = g4[22] | p4[22]&g4[6], g5[21] = g4[21] | p4[21]&g4[5], g5[20] = g4[20] | p4[20]&g4[4], g5[19] = g4[19] | p4[19]&g4[3], g5[18] = g4[18] | p4[18]&g4[2], g5[17] = g4[17] | p4[17]&g4[1], g5[16] = g4[16] | p4[16]&g4[0], g5[15] = g4[15], g5[14] = g4[14], g5[13] = g4[13], g5[12] = g4[12], g5[11] = g4[11], g5[10] = g4[10], g5[9] = g4[9], g5[8] = g4[8], g5[7] = g4[7], g5[6] = g4[6], g5[5] = g4[5], g5[4] = g4[4], g5[3] = g4[3], g5[2] = g4[2], g5[1] = g4[1], g5[0] = g4[0];
	assign p5[31] = p4[31]&p4[15], p5[30] = p4[30]&p4[14], p5[29] = p4[29]&p4[13], p5[28] = p4[28]&p4[12], p5[27] = p4[27]&p4[11], p5[26] = p4[26]&p4[10], p5[25] = p4[25]&p4[9], p5[24] = p4[24]&p4[8], p5[23] = p4[23]&p4[7], p5[22] = p4[22]&p4[6], p5[21] = p4[21]&p4[5], p5[20] = p4[20]&p4[4], p5[19] = p4[19]&p4[3], p5[18] = p4[18]&p4[2], p5[17] = p4[17]&p4[1], p5[16] = p4[16]&p4[0], p5[15] = p4[15], p5[14] = p4[14], p5[13] = p4[13], p5[12] = p4[12], p5[11] = p4[11], p5[10] = p4[10], p5[9] = p4[9], p5[8] = p4[8], p5[7] = p4[7], p5[6] = p4[6], p5[5] = p4[5], p5[4] = p4[4], p5[3] = p4[3], p5[2] = p4[2], p5[1] = p4[1], p5[0] = p4[0];



	assign c[32:1] = g5[31:0];
	assign s = p0^c[31:0];
	assign cOut = c[32];

endmodule
