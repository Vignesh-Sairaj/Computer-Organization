module Prefix_Add16(x, y, cIn, s, cOut);

	input [15:0] x, y;
	input cIn;

	output [15:0] s;
	output cOut;

	wire [15:0] g0, p0, g1, p1, g2, p2, g3, p3, g4, p4;
	wire [16:0] c;

	assign g0[15:1] = x[15:1]&y[15:1];
	assign p0[15:0] = x^y;
	assign c[0] = cIn;
	assign g0[0] = x[0]&y[0] | c[0]&(x[0] | y[0]);



	assign g1[15] = g0[15] | p0[15]&g0[14], g1[14] = g0[14] | p0[14]&g0[13], g1[13] = g0[13] | p0[13]&g0[12], g1[12] = g0[12] | p0[12]&g0[11], g1[11] = g0[11] | p0[11]&g0[10], g1[10] = g0[10] | p0[10]&g0[9], g1[9] = g0[9] | p0[9]&g0[8], g1[8] = g0[8] | p0[8]&g0[7], g1[7] = g0[7] | p0[7]&g0[6], g1[6] = g0[6] | p0[6]&g0[5], g1[5] = g0[5] | p0[5]&g0[4], g1[4] = g0[4] | p0[4]&g0[3], g1[3] = g0[3] | p0[3]&g0[2], g1[2] = g0[2] | p0[2]&g0[1], g1[1] = g0[1] | p0[1]&g0[0], g1[0] = g0[0];
	assign p1[15] = p0[15]&p0[14], p1[14] = p0[14]&p0[13], p1[13] = p0[13]&p0[12], p1[12] = p0[12]&p0[11], p1[11] = p0[11]&p0[10], p1[10] = p0[10]&p0[9], p1[9] = p0[9]&p0[8], p1[8] = p0[8]&p0[7], p1[7] = p0[7]&p0[6], p1[6] = p0[6]&p0[5], p1[5] = p0[5]&p0[4], p1[4] = p0[4]&p0[3], p1[3] = p0[3]&p0[2], p1[2] = p0[2]&p0[1], p1[1] = p0[1]&p0[0], p1[0] = p0[0];

	assign g2[15] = g1[15] | p1[15]&g1[13], g2[14] = g1[14] | p1[14]&g1[12], g2[13] = g1[13] | p1[13]&g1[11], g2[12] = g1[12] | p1[12]&g1[10], g2[11] = g1[11] | p1[11]&g1[9], g2[10] = g1[10] | p1[10]&g1[8], g2[9] = g1[9] | p1[9]&g1[7], g2[8] = g1[8] | p1[8]&g1[6], g2[7] = g1[7] | p1[7]&g1[5], g2[6] = g1[6] | p1[6]&g1[4], g2[5] = g1[5] | p1[5]&g1[3], g2[4] = g1[4] | p1[4]&g1[2], g2[3] = g1[3] | p1[3]&g1[1], g2[2] = g1[2] | p1[2]&g1[0], g2[1] = g1[1], g2[0] = g1[0];
	assign p2[15] = p1[15]&p1[13], p2[14] = p1[14]&p1[12], p2[13] = p1[13]&p1[11], p2[12] = p1[12]&p1[10], p2[11] = p1[11]&p1[9], p2[10] = p1[10]&p1[8], p2[9] = p1[9]&p1[7], p2[8] = p1[8]&p1[6], p2[7] = p1[7]&p1[5], p2[6] = p1[6]&p1[4], p2[5] = p1[5]&p1[3], p2[4] = p1[4]&p1[2], p2[3] = p1[3]&p1[1], p2[2] = p1[2]&p1[0], p2[1] = p1[1], p2[0] = p1[0];

	assign g3[15] = g2[15] | p2[15]&g2[11], g3[14] = g2[14] | p2[14]&g2[10], g3[13] = g2[13] | p2[13]&g2[9], g3[12] = g2[12] | p2[12]&g2[8], g3[11] = g2[11] | p2[11]&g2[7], g3[10] = g2[10] | p2[10]&g2[6], g3[9] = g2[9] | p2[9]&g2[5], g3[8] = g2[8] | p2[8]&g2[4], g3[7] = g2[7] | p2[7]&g2[3], g3[6] = g2[6] | p2[6]&g2[2], g3[5] = g2[5] | p2[5]&g2[1], g3[4] = g2[4] | p2[4]&g2[0], g3[3] = g2[3], g3[2] = g2[2], g3[1] = g2[1], g3[0] = g2[0];
	assign p3[15] = p2[15]&p2[11], p3[14] = p2[14]&p2[10], p3[13] = p2[13]&p2[9], p3[12] = p2[12]&p2[8], p3[11] = p2[11]&p2[7], p3[10] = p2[10]&p2[6], p3[9] = p2[9]&p2[5], p3[8] = p2[8]&p2[4], p3[7] = p2[7]&p2[3], p3[6] = p2[6]&p2[2], p3[5] = p2[5]&p2[1], p3[4] = p2[4]&p2[0], p3[3] = p2[3], p3[2] = p2[2], p3[1] = p2[1], p3[0] = p2[0];

	assign g4[15] = g3[15] | p3[15]&g3[7], g4[14] = g3[14] | p3[14]&g3[6], g4[13] = g3[13] | p3[13]&g3[5], g4[12] = g3[12] | p3[12]&g3[4], g4[11] = g3[11] | p3[11]&g3[3], g4[10] = g3[10] | p3[10]&g3[2], g4[9] = g3[9] | p3[9]&g3[1], g4[8] = g3[8] | p3[8]&g3[0], g4[7] = g3[7], g4[6] = g3[6], g4[5] = g3[5], g4[4] = g3[4], g4[3] = g3[3], g4[2] = g3[2], g4[1] = g3[1], g4[0] = g3[0];
	assign p4[15] = p3[15]&p3[7], p4[14] = p3[14]&p3[6], p4[13] = p3[13]&p3[5], p4[12] = p3[12]&p3[4], p4[11] = p3[11]&p3[3], p4[10] = p3[10]&p3[2], p4[9] = p3[9]&p3[1], p4[8] = p3[8]&p3[0], p4[7] = p3[7], p4[6] = p3[6], p4[5] = p3[5], p4[4] = p3[4], p4[3] = p3[3], p4[2] = p3[2], p4[1] = p3[1], p4[0] = p3[0];



	assign c[16:1] = g4[15:0];
	assign s = p0^c[15:0];
	assign cOut = c[16];

endmodule
